LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.all;

ENTITY L6 IS
	PORT( S :    IN STD_LOGIC_VECTOR(2 DOWNTO 0);
			E :    IN STD_LOGIC;
			F :    OUT STD_LOGIC);
END L6;

ARCHITECTURE Behavior OF L6 IS
	COMPONENT T6
	PORT ( 	I :        IN STD_LOGIC_VECTOR(7 DOWNTO 0);
			E :        IN STD_LOGIC;
			S :        IN STD_LOGIC_VECTOR(2 DOWNTO 0);
			Z :        OUT STD_LOGIC) ;
	END COMPONENT;
	
	BEGIN
		MUX: T6 PORT MAP ("11100011",E, S, F);
END Behavior;
		
	
		
			